module no2

  (input ck, //輸入外部時鐘 pin43
   output reg[6:0] s,//輸出 七段顯示器
   input [3:0] R,//輸入 偵測 row 橫列
   output reg [2:0] C);//輸出  掃描 colum 直行

  reg [13:0] t; //計數暫存器(除頻用)
  always@(posedge ck)t<=t+1;//計數 外部時鐘上緣觸發
  always@(posedge t[13])//七段掃描 自訂時鐘(t[13])上緣觸發

  case(C) //掃描 colum 直行

    3'b001:
    begin //當列輸出 第一列 High

      C<=3'b010; //下一步

      if(R==4'b0001)
        s<=7'b1111001; //1

      if(R==4'b0010)
        s<=7'b0011001; //4

      if(R==4'b0100)
        s<=7'b1111000; //7

      if(R==4'b1000)
        s<=7'b0110010; //*
    end

    3'b010:
    begin //當列輸出 第二列 High

      C<=3'b100;//下一步

      if(R==4'b0001)//判斷鍵盤行輸入 第二列High 且 第一行High 時
        s<=7'b0100100;//2

      if(R==4'b0010)//判斷鍵盤行輸入 第二列High 且 第二行High 時
        s<=7'b0010010;//5

      if(R==4'b0100)//判斷鍵盤行輸入 第二列High 且 第三行High 時
        s<=7'b0000000;//8

      if(R==4'b1000)//判斷鍵盤行輸入 第一列High 且 第三行High 時
        s<=7'b1000000;//0
    end

    default:
    begin //當列輸出 第三列 High

      C<=3'b001;//下一步

      if(R==4'b0001)//判斷鍵盤行輸入 第三列High 且 第一行High 時
        s<=7'b0110000;//3

      if(R==4'b0010)//判斷鍵盤行輸入 第三列High 且 第二行High 時
        s<=7'b0000011;//6

      if(R==4'b0100)//判斷鍵盤行輸入 第三列High 且 第三行High 時
        s<=7'b0011000;//9

      if(R==4'b1000)//判斷鍵盤行輸入 第一列High 且 第三行High 時
        s<=7'b1110000;//#
    end

  endcase
endmodule
